module complementary_filter(
  input wire clk_100mhz,
  input wire rst_in,
  input wire [15:0] gx,
  input wire [15:0] gy,
  input wire [15:0] gz,
  input wire [15:0] ax,
  input wire [15:0] ay,
  input wire [15:0] az,
)